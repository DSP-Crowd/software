-- altremote.vhd

-- Generated using ACDS version 14.0 200 at 2016.01.05.01:23:59

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altremote is
	port (
		read_param  : in  std_logic                     := '0';             --  read_param.read_param
		param       : in  std_logic_vector(2 downto 0)  := (others => '0'); --       param.param
		reconfig    : in  std_logic                     := '0';             --    reconfig.reconfig
		reset_timer : in  std_logic                     := '0';             -- reset_timer.reset_timer
		clock       : in  std_logic                     := '0';             --       clock.clk
		reset       : in  std_logic                     := '0';             --       reset.reset
		busy        : out std_logic;                                        --        busy.busy
		data_out    : out std_logic_vector(28 downto 0);                    --    data_out.data_out
		read_source : in  std_logic_vector(1 downto 0)  := (others => '0'); -- read_source.read_source
		write_param : in  std_logic                     := '0';             -- write_param.write_param
		data_in     : in  std_logic_vector(23 downto 0) := (others => '0')  --     data_in.data_in
	);
end entity altremote;

architecture rtl of altremote is
	component altremote_remote_update_0 is
		port (
			read_param  : in  std_logic                     := 'X';             -- read_param
			param       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- param
			reconfig    : in  std_logic                     := 'X';             -- reconfig
			reset_timer : in  std_logic                     := 'X';             -- reset_timer
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			busy        : out std_logic;                                        -- busy
			data_out    : out std_logic_vector(28 downto 0);                    -- data_out
			read_source : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- read_source
			write_param : in  std_logic                     := 'X';             -- write_param
			data_in     : in  std_logic_vector(23 downto 0) := (others => 'X')  -- data_in
		);
	end component altremote_remote_update_0;

begin

	remote_update_0 : component altremote_remote_update_0
		port map (
			read_param  => read_param,  --  read_param.read_param
			param       => param,       --       param.param
			reconfig    => reconfig,    --    reconfig.reconfig
			reset_timer => reset_timer, -- reset_timer.reset_timer
			clock       => clock,       --       clock.clk
			reset       => reset,       --       reset.reset
			busy        => busy,        --        busy.busy
			data_out    => data_out,    --    data_out.data_out
			read_source => read_source, -- read_source.read_source
			write_param => write_param, -- write_param.write_param
			data_in     => data_in      --     data_in.data_in
		);

end architecture rtl; -- of altremote
